library ieee;
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;


entity gh_round_perm_logic is --������������	���	�������	P	� �������������� (�������������� ������������).

port (
	after_s	: in std_logic_vector(511 downto 0);
	after_p	: out std_logic_vector(511 downto 0)
);
	end gh_round_perm_logic;
	
	--�������� ��������� ������� �� ����:
	architecture arch of gh_round_perm_logic is
	type mass_7x7_type is array (0 to 7) of std_logic_vector(7 downto 0);
	
	--�������� ���������� ������� �� ����:
	
	type mass_7x7x7_type is array (0 to 7) of mass_7x7_type;
	signal after_s_int : mass_7x7x7_type := (others => (others => (others => '0')));
	signal after_p_int : mass_7x7x7_type := (others => (others => (others => '0')));

 
begin
	--�������������� ������������� ������ �� �������� ������� � �����
 	--����������	�������	���	����,	�����	�������	������	512	�������� ������������ ���������
 	
 	fill_inputs_cycle_i: for in_i in 0 to 7 generate fill_inputs_cycle_j: for in_j in 0 to 7 generate  after_s_int(in_i)(in_j)	<= after_s((7+in_i*64+in_j*8) downto in_i*64+in_j*8);

	end generate fill_inputs_cycle_j; 
	end generate fill_inputs_cycle_i;

	--�������������� ���������� ��������� ������:
	
	rotate_cycle_i: for in_i in 0 to 7 generate rotate_cycle_j: for in_j in 0 to 7 generate after_p_int(in_j)(in_i) <= after_s_int(in_i)(in_j); 
	end generate rotate_cycle_j;
	end generate rotate_cycle_i;
	
	--�������������� ������������� ������ ��������� �� ������� � �������� ������ ��� ����, 
	--����� ������������ �� ���������� ������� ������ ������� 512-��������� ������
	
	fill_outputs_cycle_i: for in_i in 0 to 7 generate fill_outputs_cycle_j: for in_j in 0 to 7 generate after_p((7+in_i*64+in_j*8) downto in_i*64+in_j*8) <= after_p_int(in_i)(in_j);
	end generate fill_outputs_cycle_j; 
	end generate fill_outputs_cycle_i;	
end arch;

