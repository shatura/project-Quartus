module FormImp( //������� ������ � ������ FormImp
input logic clk, reset, //������������� �����
output logic [7:0]GPIO //� ������
);
logic [3:0] i; //������� ������� 4 ��� ��� ��������
				//��������� ��������
logic [15:0] X; //������� ������� 16 ��� ��� ��������
				//��������� �����������
always_ff@(posedge clk, posedge reset) //������� �������
begin
if(reset) i = 4'b0000;
else i = i + 4'b0001;
end
always_comb 	//������� ����������
begin
case(i)
4'b0000: X = 16'b0000000000000001;
4'b0001: X = 16'b0000000000000010;
4'b0010: X = 16'b0000000000000100;
4'b0011: X = 16'b0000000000001000;
4'b0100: X = 16'b0000000000010000;
4'b0101: X = 16'b0000000000100000;
4'b0110: X = 16'b0000000001000000;
4'b0111: X = 16'b0000000010000000;
4'b1000: X = 16'b0000000100000000;
4'b1001: X = 16'b0000001000000000;
4'b1010: X = 16'b0000010000000000;
4'b1011: X = 16'b0000100000000000;
4'b1100: X = 16'b0001000000000000;
4'b1101: X = 16'b0010000000000000;
4'b1110: X = 16'b0100000000000000;
4'b1111: X = 16'b1000000000000000;
endcase
end
always_ff@(posedge X[0], posedge X[8]) //����� �������� ����������
										//� 0-��
begin 									//� 8-�� ������ �����������
if (X[0]) GPIO[0] <= 1; 		//���������
else if (X[8]) GPIO[0] <= 0; 	//�����
end
always_ff@(posedge X[1], posedge X[9]) //����� �������� ����������
										//� 1-��
begin 									//� 9-�� ������ �����������
if (X[1]) GPIO[1] <= 1; //���������
else if (X[9]) GPIO[1] <= 0; //�����
end
always_ff@(posedge X[2], posedge X[10]) //����� �������� ����������
										//� 2-�� �10-��
begin 									//������ �����������
if (X[2]) GPIO[2] <= 1; //���������
else if (X[10]) GPIO[2] <= 0; //�����
end
always_ff@(posedge X[3], posedge X[11]) //����� �������� ����������
										//� 3-�� � 11-��
begin									 //������ �����������
if (X[3]) GPIO[3] <= 1; //���������
else if (X[11]) GPIO[3] <= 0; //�����
end
always_ff@(posedge X[4], posedge X[12]) //����� �������� ����������
										//� 4-�� � 12-��
begin 									// ������ �����������
if (X[4]) GPIO[4] <= 1; //���������
else if (X[12]) GPIO[4] <= 0; //�����
end
always_ff@(posedge X[5], posedge X[13]) //����� �������� ����������
										//� 5-�� � 13-��
begin 									// ������ �����������
if (X[5]) GPIO[5] <= 1; //���������
else if (X[13]) GPIO[5] <= 0; //�����
end
always_ff@(posedge X[6], posedge X[14]) //����� �������� ����������
										//� 6-�� � 14-��
begin 									//������ �����������
if (X[6]) GPIO[6] <= 1; //���������
else if (X[14]) GPIO[6] <= 0; //�����
end
always_ff@(posedge X[7], posedge X[15]) //����� �������� ����������
										//� 7-�� � 15-��
begin 									// ������ �����������
if (X[7]) GPIO[7] <= 1; //���������
else if (X[15]) GPIO[7] <= 0; //�����
end
endmodule //����� ������